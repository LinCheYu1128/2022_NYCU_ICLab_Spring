module div_3_12b(
	input [11:0]in,
	output reg[10:0]out
);
	always@(in)
		case(in)
			12'b111111101100:out = 10'b1111111010;        //-20/3=-6
			12'b111111101101:out = 10'b1111111010;        //-19/3=-6
			12'b111111101110:out = 10'b1111111010;        //-18/3=-6
			12'b111111101111:out = 10'b1111111011;        //-17/3=-5
			12'b111111110000:out = 10'b1111111011;        //-16/3=-5
			12'b111111110001:out = 10'b1111111011;        //-15/3=-5
			12'b111111110010:out = 10'b1111111100;        //-14/3=-4
			12'b111111110011:out = 10'b1111111100;        //-13/3=-4
			12'b111111110100:out = 10'b1111111100;        //-12/3=-4
			12'b111111110101:out = 10'b1111111101;        //-11/3=-3
			12'b111111110110:out = 10'b1111111101;        //-10/3=-3
			12'b111111110111:out = 10'b1111111101;        //-9/3=-3
			12'b111111111000:out = 10'b1111111110;        //-8/3=-2
			12'b111111111001:out = 10'b1111111110;        //-7/3=-2
			12'b111111111010:out = 10'b1111111110;        //-6/3=-2
			12'b111111111011:out = 10'b1111111111;        //-5/3=-1
			12'b111111111100:out = 10'b1111111111;        //-4/3=-1
			12'b111111111101:out = 10'b1111111111;        //-3/3=-1
			12'b111111111110:out = 10'b0000000000;        //-2/3=0
			12'b111111111111:out = 10'b0000000000;        //-1/3=0
			12'b000000000000:out = 10'b0000000000;        //0/3=0
			12'b000000000001:out = 10'b0000000000;        //1/3=0
			12'b000000000010:out = 10'b0000000000;        //2/3=0
			12'b000000000011:out = 10'b0000000001;        //3/3=1
			12'b000000000100:out = 10'b0000000001;        //4/3=1
			12'b000000000101:out = 10'b0000000001;        //5/3=1
			12'b000000000110:out = 10'b0000000010;        //6/3=2
			12'b000000000111:out = 10'b0000000010;        //7/3=2
			12'b000000001000:out = 10'b0000000010;        //8/3=2
			12'b000000001001:out = 10'b0000000011;        //9/3=3
			12'b000000001010:out = 10'b0000000011;        //10/3=3
			12'b000000001011:out = 10'b0000000011;        //11/3=3
			12'b000000001100:out = 10'b0000000100;        //12/3=4
			12'b000000001101:out = 10'b0000000100;        //13/3=4
			12'b000000001110:out = 10'b0000000100;        //14/3=4
			12'b000000001111:out = 10'b0000000101;        //15/3=5
			12'b000000010000:out = 10'b0000000101;        //16/3=5
			12'b000000010001:out = 10'b0000000101;        //17/3=5
			12'b000000010010:out = 10'b0000000110;        //18/3=6
			12'b000000010011:out = 10'b0000000110;        //19/3=6
			12'b000000010100:out = 10'b0000000110;        //20/3=6
			12'b000000010101:out = 10'b0000000111;        //21/3=7
			12'b000000010110:out = 10'b0000000111;        //22/3=7
			12'b000000010111:out = 10'b0000000111;        //23/3=7
			12'b000000011000:out = 10'b0000001000;        //24/3=8
			12'b000000011001:out = 10'b0000001000;        //25/3=8
			12'b000000011010:out = 10'b0000001000;        //26/3=8
			12'b000000011011:out = 10'b0000001001;        //27/3=9
			12'b000000011100:out = 10'b0000001001;        //28/3=9
			12'b000000011101:out = 10'b0000001001;        //29/3=9
			12'b000000011110:out = 10'b0000001010;        //30/3=10
			12'b000000011111:out = 10'b0000001010;        //31/3=10
			12'b000000100000:out = 10'b0000001010;        //32/3=10
			12'b000000100001:out = 10'b0000001011;        //33/3=11
			12'b000000100010:out = 10'b0000001011;        //34/3=11
			12'b000000100011:out = 10'b0000001011;        //35/3=11
			12'b000000100100:out = 10'b0000001100;        //36/3=12
			12'b000000100101:out = 10'b0000001100;        //37/3=12
			12'b000000100110:out = 10'b0000001100;        //38/3=12
			12'b000000100111:out = 10'b0000001101;        //39/3=13
			12'b000000101000:out = 10'b0000001101;        //40/3=13
			12'b000000101001:out = 10'b0000001101;        //41/3=13
			12'b000000101010:out = 10'b0000001110;        //42/3=14
			12'b000000101011:out = 10'b0000001110;        //43/3=14
			12'b000000101100:out = 10'b0000001110;        //44/3=14
			12'b000000101101:out = 10'b0000001111;        //45/3=15
			12'b000000101110:out = 10'b0000001111;        //46/3=15
			12'b000000101111:out = 10'b0000001111;        //47/3=15
			12'b000000110000:out = 10'b0000010000;        //48/3=16
			12'b000000110001:out = 10'b0000010000;        //49/3=16
			12'b000000110010:out = 10'b0000010000;        //50/3=16
			12'b000000110011:out = 10'b0000010001;        //51/3=17
			12'b000000110100:out = 10'b0000010001;        //52/3=17
			12'b000000110101:out = 10'b0000010001;        //53/3=17
			12'b000000110110:out = 10'b0000010010;        //54/3=18
			12'b000000110111:out = 10'b0000010010;        //55/3=18
			12'b000000111000:out = 10'b0000010010;        //56/3=18
			12'b000000111001:out = 10'b0000010011;        //57/3=19
			12'b000000111010:out = 10'b0000010011;        //58/3=19
			12'b000000111011:out = 10'b0000010011;        //59/3=19
			12'b000000111100:out = 10'b0000010100;        //60/3=20
			12'b000000111101:out = 10'b0000010100;        //61/3=20
			12'b000000111110:out = 10'b0000010100;        //62/3=20
			12'b000000111111:out = 10'b0000010101;        //63/3=21
			12'b000001000000:out = 10'b0000010101;        //64/3=21
			12'b000001000001:out = 10'b0000010101;        //65/3=21
			12'b000001000010:out = 10'b0000010110;        //66/3=22
			12'b000001000011:out = 10'b0000010110;        //67/3=22
			12'b000001000100:out = 10'b0000010110;        //68/3=22
			12'b000001000101:out = 10'b0000010111;        //69/3=23
			12'b000001000110:out = 10'b0000010111;        //70/3=23
			12'b000001000111:out = 10'b0000010111;        //71/3=23
			12'b000001001000:out = 10'b0000011000;        //72/3=24
			12'b000001001001:out = 10'b0000011000;        //73/3=24
			12'b000001001010:out = 10'b0000011000;        //74/3=24
			12'b000001001011:out = 10'b0000011001;        //75/3=25
			12'b000001001100:out = 10'b0000011001;        //76/3=25
			12'b000001001101:out = 10'b0000011001;        //77/3=25
			12'b000001001110:out = 10'b0000011010;        //78/3=26
			12'b000001001111:out = 10'b0000011010;        //79/3=26
			12'b000001010000:out = 10'b0000011010;        //80/3=26
			12'b000001010001:out = 10'b0000011011;        //81/3=27
			12'b000001010010:out = 10'b0000011011;        //82/3=27
			12'b000001010011:out = 10'b0000011011;        //83/3=27
			12'b000001010100:out = 10'b0000011100;        //84/3=28
			12'b000001010101:out = 10'b0000011100;        //85/3=28
			12'b000001010110:out = 10'b0000011100;        //86/3=28
			12'b000001010111:out = 10'b0000011101;        //87/3=29
			12'b000001011000:out = 10'b0000011101;        //88/3=29
			12'b000001011001:out = 10'b0000011101;        //89/3=29
			12'b000001011010:out = 10'b0000011110;        //90/3=30
			12'b000001011011:out = 10'b0000011110;        //91/3=30
			12'b000001011100:out = 10'b0000011110;        //92/3=30
			12'b000001011101:out = 10'b0000011111;        //93/3=31
			12'b000001011110:out = 10'b0000011111;        //94/3=31
			12'b000001011111:out = 10'b0000011111;        //95/3=31
			12'b000001100000:out = 10'b0000100000;        //96/3=32
			12'b000001100001:out = 10'b0000100000;        //97/3=32
			12'b000001100010:out = 10'b0000100000;        //98/3=32
			12'b000001100011:out = 10'b0000100001;        //99/3=33
			12'b000001100100:out = 10'b0000100001;        //100/3=33
			12'b000001100101:out = 10'b0000100001;        //101/3=33
			12'b000001100110:out = 10'b0000100010;        //102/3=34
			12'b000001100111:out = 10'b0000100010;        //103/3=34
			12'b000001101000:out = 10'b0000100010;        //104/3=34
			12'b000001101001:out = 10'b0000100011;        //105/3=35
			12'b000001101010:out = 10'b0000100011;        //106/3=35
			12'b000001101011:out = 10'b0000100011;        //107/3=35
			12'b000001101100:out = 10'b0000100100;        //108/3=36
			12'b000001101101:out = 10'b0000100100;        //109/3=36
			12'b000001101110:out = 10'b0000100100;        //110/3=36
			12'b000001101111:out = 10'b0000100101;        //111/3=37
			12'b000001110000:out = 10'b0000100101;        //112/3=37
			12'b000001110001:out = 10'b0000100101;        //113/3=37
			12'b000001110010:out = 10'b0000100110;        //114/3=38
			12'b000001110011:out = 10'b0000100110;        //115/3=38
			12'b000001110100:out = 10'b0000100110;        //116/3=38
			12'b000001110101:out = 10'b0000100111;        //117/3=39
			12'b000001110110:out = 10'b0000100111;        //118/3=39
			12'b000001110111:out = 10'b0000100111;        //119/3=39
			12'b000001111000:out = 10'b0000101000;        //120/3=40
			12'b000001111001:out = 10'b0000101000;        //121/3=40
			12'b000001111010:out = 10'b0000101000;        //122/3=40
			12'b000001111011:out = 10'b0000101001;        //123/3=41
			12'b000001111100:out = 10'b0000101001;        //124/3=41
			12'b000001111101:out = 10'b0000101001;        //125/3=41
			12'b000001111110:out = 10'b0000101010;        //126/3=42
			12'b000001111111:out = 10'b0000101010;        //127/3=42
			12'b000010000000:out = 10'b0000101010;        //128/3=42
			12'b000010000001:out = 10'b0000101011;        //129/3=43
			12'b000010000010:out = 10'b0000101011;        //130/3=43
			12'b000010000011:out = 10'b0000101011;        //131/3=43
			12'b000010000100:out = 10'b0000101100;        //132/3=44
			12'b000010000101:out = 10'b0000101100;        //133/3=44
			12'b000010000110:out = 10'b0000101100;        //134/3=44
			12'b000010000111:out = 10'b0000101101;        //135/3=45
			12'b000010001000:out = 10'b0000101101;        //136/3=45
			12'b000010001001:out = 10'b0000101101;        //137/3=45
			12'b000010001010:out = 10'b0000101110;        //138/3=46
			12'b000010001011:out = 10'b0000101110;        //139/3=46
			12'b000010001100:out = 10'b0000101110;        //140/3=46
			12'b000010001101:out = 10'b0000101111;        //141/3=47
			12'b000010001110:out = 10'b0000101111;        //142/3=47
			12'b000010001111:out = 10'b0000101111;        //143/3=47
			12'b000010010000:out = 10'b0000110000;        //144/3=48
			12'b000010010001:out = 10'b0000110000;        //145/3=48
			12'b000010010010:out = 10'b0000110000;        //146/3=48
			12'b000010010011:out = 10'b0000110001;        //147/3=49
			12'b000010010100:out = 10'b0000110001;        //148/3=49
			12'b000010010101:out = 10'b0000110001;        //149/3=49
			12'b000010010110:out = 10'b0000110010;        //150/3=50
			12'b000010010111:out = 10'b0000110010;        //151/3=50
			12'b000010011000:out = 10'b0000110010;        //152/3=50
			12'b000010011001:out = 10'b0000110011;        //153/3=51
			12'b000010011010:out = 10'b0000110011;        //154/3=51
			12'b000010011011:out = 10'b0000110011;        //155/3=51
			12'b000010011100:out = 10'b0000110100;        //156/3=52
			12'b000010011101:out = 10'b0000110100;        //157/3=52
			12'b000010011110:out = 10'b0000110100;        //158/3=52
			12'b000010011111:out = 10'b0000110101;        //159/3=53
			12'b000010100000:out = 10'b0000110101;        //160/3=53
			12'b000010100001:out = 10'b0000110101;        //161/3=53
			12'b000010100010:out = 10'b0000110110;        //162/3=54
			12'b000010100011:out = 10'b0000110110;        //163/3=54
			12'b000010100100:out = 10'b0000110110;        //164/3=54
			12'b000010100101:out = 10'b0000110111;        //165/3=55
			12'b000010100110:out = 10'b0000110111;        //166/3=55
			12'b000010100111:out = 10'b0000110111;        //167/3=55
			12'b000010101000:out = 10'b0000111000;        //168/3=56
			12'b000010101001:out = 10'b0000111000;        //169/3=56
			12'b000010101010:out = 10'b0000111000;        //170/3=56
			12'b000010101011:out = 10'b0000111001;        //171/3=57
			12'b000010101100:out = 10'b0000111001;        //172/3=57
			12'b000010101101:out = 10'b0000111001;        //173/3=57
			12'b000010101110:out = 10'b0000111010;        //174/3=58
			12'b000010101111:out = 10'b0000111010;        //175/3=58
			12'b000010110000:out = 10'b0000111010;        //176/3=58
			12'b000010110001:out = 10'b0000111011;        //177/3=59
			12'b000010110010:out = 10'b0000111011;        //178/3=59
			12'b000010110011:out = 10'b0000111011;        //179/3=59
			12'b000010110100:out = 10'b0000111100;        //180/3=60
			12'b000010110101:out = 10'b0000111100;        //181/3=60
			12'b000010110110:out = 10'b0000111100;        //182/3=60
			12'b000010110111:out = 10'b0000111101;        //183/3=61
			12'b000010111000:out = 10'b0000111101;        //184/3=61
			12'b000010111001:out = 10'b0000111101;        //185/3=61
			12'b000010111010:out = 10'b0000111110;        //186/3=62
			12'b000010111011:out = 10'b0000111110;        //187/3=62
			12'b000010111100:out = 10'b0000111110;        //188/3=62
			12'b000010111101:out = 10'b0000111111;        //189/3=63
			12'b000010111110:out = 10'b0000111111;        //190/3=63
			12'b000010111111:out = 10'b0000111111;        //191/3=63
			12'b000011000000:out = 10'b0001000000;        //192/3=64
			12'b000011000001:out = 10'b0001000000;        //193/3=64
			12'b000011000010:out = 10'b0001000000;        //194/3=64
			12'b000011000011:out = 10'b0001000001;        //195/3=65
			12'b000011000100:out = 10'b0001000001;        //196/3=65
			12'b000011000101:out = 10'b0001000001;        //197/3=65
			12'b000011000110:out = 10'b0001000010;        //198/3=66
			12'b000011000111:out = 10'b0001000010;        //199/3=66
			12'b000011001000:out = 10'b0001000010;        //200/3=66
			12'b000011001001:out = 10'b0001000011;        //201/3=67
			12'b000011001010:out = 10'b0001000011;        //202/3=67
			12'b000011001011:out = 10'b0001000011;        //203/3=67
			12'b000011001100:out = 10'b0001000100;        //204/3=68
			12'b000011001101:out = 10'b0001000100;        //205/3=68
			12'b000011001110:out = 10'b0001000100;        //206/3=68
			12'b000011001111:out = 10'b0001000101;        //207/3=69
			12'b000011010000:out = 10'b0001000101;        //208/3=69
			12'b000011010001:out = 10'b0001000101;        //209/3=69
			12'b000011010010:out = 10'b0001000110;        //210/3=70
			12'b000011010011:out = 10'b0001000110;        //211/3=70
			12'b000011010100:out = 10'b0001000110;        //212/3=70
			12'b000011010101:out = 10'b0001000111;        //213/3=71
			12'b000011010110:out = 10'b0001000111;        //214/3=71
			12'b000011010111:out = 10'b0001000111;        //215/3=71
			12'b000011011000:out = 10'b0001001000;        //216/3=72
			12'b000011011001:out = 10'b0001001000;        //217/3=72
			12'b000011011010:out = 10'b0001001000;        //218/3=72
			12'b000011011011:out = 10'b0001001001;        //219/3=73
			12'b000011011100:out = 10'b0001001001;        //220/3=73
			12'b000011011101:out = 10'b0001001001;        //221/3=73
			12'b000011011110:out = 10'b0001001010;        //222/3=74
			12'b000011011111:out = 10'b0001001010;        //223/3=74
			12'b000011100000:out = 10'b0001001010;        //224/3=74
			12'b000011100001:out = 10'b0001001011;        //225/3=75
			12'b000011100010:out = 10'b0001001011;        //226/3=75
			12'b000011100011:out = 10'b0001001011;        //227/3=75
			12'b000011100100:out = 10'b0001001100;        //228/3=76
			12'b000011100101:out = 10'b0001001100;        //229/3=76
			12'b000011100110:out = 10'b0001001100;        //230/3=76
			12'b000011100111:out = 10'b0001001101;        //231/3=77
			12'b000011101000:out = 10'b0001001101;        //232/3=77
			12'b000011101001:out = 10'b0001001101;        //233/3=77
			12'b000011101010:out = 10'b0001001110;        //234/3=78
			12'b000011101011:out = 10'b0001001110;        //235/3=78
			12'b000011101100:out = 10'b0001001110;        //236/3=78
			12'b000011101101:out = 10'b0001001111;        //237/3=79
			12'b000011101110:out = 10'b0001001111;        //238/3=79
			12'b000011101111:out = 10'b0001001111;        //239/3=79
			12'b000011110000:out = 10'b0001010000;        //240/3=80
			12'b000011110001:out = 10'b0001010000;        //241/3=80
			12'b000011110010:out = 10'b0001010000;        //242/3=80
			12'b000011110011:out = 10'b0001010001;        //243/3=81
			12'b000011110100:out = 10'b0001010001;        //244/3=81
			12'b000011110101:out = 10'b0001010001;        //245/3=81
			12'b000011110110:out = 10'b0001010010;        //246/3=82
			12'b000011110111:out = 10'b0001010010;        //247/3=82
			12'b000011111000:out = 10'b0001010010;        //248/3=82
			12'b000011111001:out = 10'b0001010011;        //249/3=83
			12'b000011111010:out = 10'b0001010011;        //250/3=83
			12'b000011111011:out = 10'b0001010011;        //251/3=83
			12'b000011111100:out = 10'b0001010100;        //252/3=84
			12'b000011111101:out = 10'b0001010100;        //253/3=84
			12'b000011111110:out = 10'b0001010100;        //254/3=84
			12'b000011111111:out = 10'b0001010101;        //255/3=85
			12'b000100000000:out = 10'b0001010101;        //256/3=85
			12'b000100000001:out = 10'b0001010101;        //257/3=85
			12'b000100000010:out = 10'b0001010110;        //258/3=86
			12'b000100000011:out = 10'b0001010110;        //259/3=86
			12'b000100000100:out = 10'b0001010110;        //260/3=86
			12'b000100000101:out = 10'b0001010111;        //261/3=87
			12'b000100000110:out = 10'b0001010111;        //262/3=87
			12'b000100000111:out = 10'b0001010111;        //263/3=87
			12'b000100001000:out = 10'b0001011000;        //264/3=88
			12'b000100001001:out = 10'b0001011000;        //265/3=88
			12'b000100001010:out = 10'b0001011000;        //266/3=88
			12'b000100001011:out = 10'b0001011001;        //267/3=89
			12'b000100001100:out = 10'b0001011001;        //268/3=89
			12'b000100001101:out = 10'b0001011001;        //269/3=89
			12'b000100001110:out = 10'b0001011010;        //270/3=90
			12'b000100001111:out = 10'b0001011010;        //271/3=90
			12'b000100010000:out = 10'b0001011010;        //272/3=90
			12'b000100010001:out = 10'b0001011011;        //273/3=91
			12'b000100010010:out = 10'b0001011011;        //274/3=91
			12'b000100010011:out = 10'b0001011011;        //275/3=91
			12'b000100010100:out = 10'b0001011100;        //276/3=92
			12'b000100010101:out = 10'b0001011100;        //277/3=92
			12'b000100010110:out = 10'b0001011100;        //278/3=92
			12'b000100010111:out = 10'b0001011101;        //279/3=93
			12'b000100011000:out = 10'b0001011101;        //280/3=93
			12'b000100011001:out = 10'b0001011101;        //281/3=93
			12'b000100011010:out = 10'b0001011110;        //282/3=94
			12'b000100011011:out = 10'b0001011110;        //283/3=94
			12'b000100011100:out = 10'b0001011110;        //284/3=94
			12'b000100011101:out = 10'b0001011111;        //285/3=95
			12'b000100011110:out = 10'b0001011111;        //286/3=95
			12'b000100011111:out = 10'b0001011111;        //287/3=95
			12'b000100100000:out = 10'b0001100000;        //288/3=96
			12'b000100100001:out = 10'b0001100000;        //289/3=96
			12'b000100100010:out = 10'b0001100000;        //290/3=96
			12'b000100100011:out = 10'b0001100001;        //291/3=97
			12'b000100100100:out = 10'b0001100001;        //292/3=97
			12'b000100100101:out = 10'b0001100001;        //293/3=97
			12'b000100100110:out = 10'b0001100010;        //294/3=98
			12'b000100100111:out = 10'b0001100010;        //295/3=98
			12'b000100101000:out = 10'b0001100010;        //296/3=98
			12'b000100101001:out = 10'b0001100011;        //297/3=99
			12'b000100101010:out = 10'b0001100011;        //298/3=99
			12'b000100101011:out = 10'b0001100011;        //299/3=99
			12'b000100101100:out = 10'b0001100100;        //300/3=100
			12'b000100101101:out = 10'b0001100100;        //301/3=100
			12'b000100101110:out = 10'b0001100100;        //302/3=100
			12'b000100101111:out = 10'b0001100101;        //303/3=101
			12'b000100110000:out = 10'b0001100101;        //304/3=101
			12'b000100110001:out = 10'b0001100101;        //305/3=101
			12'b000100110010:out = 10'b0001100110;        //306/3=102
			12'b000100110011:out = 10'b0001100110;        //307/3=102
			12'b000100110100:out = 10'b0001100110;        //308/3=102
			12'b000100110101:out = 10'b0001100111;        //309/3=103
			12'b000100110110:out = 10'b0001100111;        //310/3=103
			12'b000100110111:out = 10'b0001100111;        //311/3=103
			12'b000100111000:out = 10'b0001101000;        //312/3=104
			12'b000100111001:out = 10'b0001101000;        //313/3=104
			12'b000100111010:out = 10'b0001101000;        //314/3=104
			12'b000100111011:out = 10'b0001101001;        //315/3=105
			12'b000100111100:out = 10'b0001101001;        //316/3=105
			12'b000100111101:out = 10'b0001101001;        //317/3=105
			12'b000100111110:out = 10'b0001101010;        //318/3=106
			12'b000100111111:out = 10'b0001101010;        //319/3=106
			12'b000101000000:out = 10'b0001101010;        //320/3=106
			12'b000101000001:out = 10'b0001101011;        //321/3=107
			12'b000101000010:out = 10'b0001101011;        //322/3=107
			12'b000101000011:out = 10'b0001101011;        //323/3=107
			12'b000101000100:out = 10'b0001101100;        //324/3=108
			12'b000101000101:out = 10'b0001101100;        //325/3=108
			12'b000101000110:out = 10'b0001101100;        //326/3=108
			12'b000101000111:out = 10'b0001101101;        //327/3=109
			12'b000101001000:out = 10'b0001101101;        //328/3=109
			12'b000101001001:out = 10'b0001101101;        //329/3=109
			12'b000101001010:out = 10'b0001101110;        //330/3=110
			12'b000101001011:out = 10'b0001101110;        //331/3=110
			12'b000101001100:out = 10'b0001101110;        //332/3=110
			12'b000101001101:out = 10'b0001101111;        //333/3=111
			12'b000101001110:out = 10'b0001101111;        //334/3=111
			12'b000101001111:out = 10'b0001101111;        //335/3=111
			12'b000101010000:out = 10'b0001110000;        //336/3=112
			12'b000101010001:out = 10'b0001110000;        //337/3=112
			12'b000101010010:out = 10'b0001110000;        //338/3=112
			12'b000101010011:out = 10'b0001110001;        //339/3=113
			12'b000101010100:out = 10'b0001110001;        //340/3=113
			12'b000101010101:out = 10'b0001110001;        //341/3=113
			12'b000101010110:out = 10'b0001110010;        //342/3=114
			12'b000101010111:out = 10'b0001110010;        //343/3=114
			12'b000101011000:out = 10'b0001110010;        //344/3=114
			12'b000101011001:out = 10'b0001110011;        //345/3=115
			12'b000101011010:out = 10'b0001110011;        //346/3=115
			12'b000101011011:out = 10'b0001110011;        //347/3=115
			12'b000101011100:out = 10'b0001110100;        //348/3=116
			12'b000101011101:out = 10'b0001110100;        //349/3=116
			12'b000101011110:out = 10'b0001110100;        //350/3=116
			12'b000101011111:out = 10'b0001110101;        //351/3=117
			12'b000101100000:out = 10'b0001110101;        //352/3=117
			12'b000101100001:out = 10'b0001110101;        //353/3=117
			12'b000101100010:out = 10'b0001110110;        //354/3=118
			12'b000101100011:out = 10'b0001110110;        //355/3=118
			12'b000101100100:out = 10'b0001110110;        //356/3=118
			12'b000101100101:out = 10'b0001110111;        //357/3=119
			12'b000101100110:out = 10'b0001110111;        //358/3=119
			12'b000101100111:out = 10'b0001110111;        //359/3=119
			12'b000101101000:out = 10'b0001111000;        //360/3=120
			12'b000101101001:out = 10'b0001111000;        //361/3=120
			12'b000101101010:out = 10'b0001111000;        //362/3=120
			12'b000101101011:out = 10'b0001111001;        //363/3=121
			12'b000101101100:out = 10'b0001111001;        //364/3=121
			12'b000101101101:out = 10'b0001111001;        //365/3=121
			12'b000101101110:out = 10'b0001111010;        //366/3=122
			12'b000101101111:out = 10'b0001111010;        //367/3=122
			12'b000101110000:out = 10'b0001111010;        //368/3=122
			12'b000101110001:out = 10'b0001111011;        //369/3=123
			12'b000101110010:out = 10'b0001111011;        //370/3=123
			12'b000101110011:out = 10'b0001111011;        //371/3=123
			12'b000101110100:out = 10'b0001111100;        //372/3=124
			12'b000101110101:out = 10'b0001111100;        //373/3=124
			12'b000101110110:out = 10'b0001111100;        //374/3=124
			12'b000101110111:out = 10'b0001111101;        //375/3=125
			12'b000101111000:out = 10'b0001111101;        //376/3=125
			12'b000101111001:out = 10'b0001111101;        //377/3=125
			12'b000101111010:out = 10'b0001111110;        //378/3=126
			12'b000101111011:out = 10'b0001111110;        //379/3=126
			12'b000101111100:out = 10'b0001111110;        //380/3=126
			12'b000101111101:out = 10'b0001111111;        //381/3=127
			12'b000101111110:out = 10'b0001111111;        //382/3=127
			12'b000101111111:out = 10'b0001111111;        //383/3=127
			12'b000110000000:out = 10'b0010000000;        //384/3=128
			12'b000110000001:out = 10'b0010000000;        //385/3=128
			12'b000110000010:out = 10'b0010000000;        //386/3=128
			12'b000110000011:out = 10'b0010000001;        //387/3=129
			12'b000110000100:out = 10'b0010000001;        //388/3=129
			12'b000110000101:out = 10'b0010000001;        //389/3=129
			12'b000110000110:out = 10'b0010000010;        //390/3=130
			12'b000110000111:out = 10'b0010000010;        //391/3=130
			12'b000110001000:out = 10'b0010000010;        //392/3=130
			12'b000110001001:out = 10'b0010000011;        //393/3=131
			12'b000110001010:out = 10'b0010000011;        //394/3=131
			12'b000110001011:out = 10'b0010000011;        //395/3=131
			12'b000110001100:out = 10'b0010000100;        //396/3=132
			12'b000110001101:out = 10'b0010000100;        //397/3=132
			12'b000110001110:out = 10'b0010000100;        //398/3=132
			12'b000110001111:out = 10'b0010000101;        //399/3=133
			12'b000110010000:out = 10'b0010000101;        //400/3=133
			12'b000110010001:out = 10'b0010000101;        //401/3=133
			12'b000110010010:out = 10'b0010000110;        //402/3=134
			12'b000110010011:out = 10'b0010000110;        //403/3=134
			12'b000110010100:out = 10'b0010000110;        //404/3=134
			12'b000110010101:out = 10'b0010000111;        //405/3=135
			12'b000110010110:out = 10'b0010000111;        //406/3=135
			12'b000110010111:out = 10'b0010000111;        //407/3=135
			12'b000110011000:out = 10'b0010001000;        //408/3=136
			12'b000110011001:out = 10'b0010001000;        //409/3=136
			12'b000110011010:out = 10'b0010001000;        //410/3=136
			12'b000110011011:out = 10'b0010001001;        //411/3=137
			12'b000110011100:out = 10'b0010001001;        //412/3=137
			12'b000110011101:out = 10'b0010001001;        //413/3=137
			12'b000110011110:out = 10'b0010001010;        //414/3=138
			12'b000110011111:out = 10'b0010001010;        //415/3=138
			12'b000110100000:out = 10'b0010001010;        //416/3=138
			12'b000110100001:out = 10'b0010001011;        //417/3=139
			12'b000110100010:out = 10'b0010001011;        //418/3=139
			12'b000110100011:out = 10'b0010001011;        //419/3=139
			12'b000110100100:out = 10'b0010001100;        //420/3=140
			12'b000110100101:out = 10'b0010001100;        //421/3=140
			12'b000110100110:out = 10'b0010001100;        //422/3=140
			12'b000110100111:out = 10'b0010001101;        //423/3=141
			12'b000110101000:out = 10'b0010001101;        //424/3=141
			12'b000110101001:out = 10'b0010001101;        //425/3=141
			12'b000110101010:out = 10'b0010001110;        //426/3=142
			12'b000110101011:out = 10'b0010001110;        //427/3=142
			12'b000110101100:out = 10'b0010001110;        //428/3=142
			12'b000110101101:out = 10'b0010001111;        //429/3=143
			12'b000110101110:out = 10'b0010001111;        //430/3=143
			12'b000110101111:out = 10'b0010001111;        //431/3=143
			12'b000110110000:out = 10'b0010010000;        //432/3=144
			12'b000110110001:out = 10'b0010010000;        //433/3=144
			12'b000110110010:out = 10'b0010010000;        //434/3=144
			12'b000110110011:out = 10'b0010010001;        //435/3=145
			12'b000110110100:out = 10'b0010010001;        //436/3=145
			12'b000110110101:out = 10'b0010010001;        //437/3=145
			12'b000110110110:out = 10'b0010010010;        //438/3=146
			12'b000110110111:out = 10'b0010010010;        //439/3=146
			12'b000110111000:out = 10'b0010010010;        //440/3=146
			12'b000110111001:out = 10'b0010010011;        //441/3=147
			12'b000110111010:out = 10'b0010010011;        //442/3=147
			12'b000110111011:out = 10'b0010010011;        //443/3=147
			12'b000110111100:out = 10'b0010010100;        //444/3=148
			12'b000110111101:out = 10'b0010010100;        //445/3=148
			12'b000110111110:out = 10'b0010010100;        //446/3=148
			12'b000110111111:out = 10'b0010010101;        //447/3=149
			12'b000111000000:out = 10'b0010010101;        //448/3=149
			12'b000111000001:out = 10'b0010010101;        //449/3=149
			12'b000111000010:out = 10'b0010010110;        //450/3=150
			12'b000111000011:out = 10'b0010010110;        //451/3=150
			12'b000111000100:out = 10'b0010010110;        //452/3=150
			12'b000111000101:out = 10'b0010010111;        //453/3=151
			12'b000111000110:out = 10'b0010010111;        //454/3=151
			12'b000111000111:out = 10'b0010010111;        //455/3=151
			12'b000111001000:out = 10'b0010011000;        //456/3=152
			12'b000111001001:out = 10'b0010011000;        //457/3=152
			12'b000111001010:out = 10'b0010011000;        //458/3=152
			12'b000111001011:out = 10'b0010011001;        //459/3=153
			12'b000111001100:out = 10'b0010011001;        //460/3=153
			12'b000111001101:out = 10'b0010011001;        //461/3=153
			12'b000111001110:out = 10'b0010011010;        //462/3=154
			12'b000111001111:out = 10'b0010011010;        //463/3=154
			12'b000111010000:out = 10'b0010011010;        //464/3=154
			12'b000111010001:out = 10'b0010011011;        //465/3=155
			12'b000111010010:out = 10'b0010011011;        //466/3=155
			12'b000111010011:out = 10'b0010011011;        //467/3=155
			12'b000111010100:out = 10'b0010011100;        //468/3=156
			12'b000111010101:out = 10'b0010011100;        //469/3=156
			12'b000111010110:out = 10'b0010011100;        //470/3=156
			12'b000111010111:out = 10'b0010011101;        //471/3=157
			12'b000111011000:out = 10'b0010011101;        //472/3=157
			12'b000111011001:out = 10'b0010011101;        //473/3=157
			12'b000111011010:out = 10'b0010011110;        //474/3=158
			12'b000111011011:out = 10'b0010011110;        //475/3=158
			12'b000111011100:out = 10'b0010011110;        //476/3=158
			12'b000111011101:out = 10'b0010011111;        //477/3=159
			12'b000111011110:out = 10'b0010011111;        //478/3=159
			12'b000111011111:out = 10'b0010011111;        //479/3=159
			12'b000111100000:out = 10'b0010100000;        //480/3=160
			12'b000111100001:out = 10'b0010100000;        //481/3=160
			12'b000111100010:out = 10'b0010100000;        //482/3=160
			12'b000111100011:out = 10'b0010100001;        //483/3=161
			12'b000111100100:out = 10'b0010100001;        //484/3=161
			12'b000111100101:out = 10'b0010100001;        //485/3=161
			12'b000111100110:out = 10'b0010100010;        //486/3=162
			12'b000111100111:out = 10'b0010100010;        //487/3=162
			12'b000111101000:out = 10'b0010100010;        //488/3=162
			12'b000111101001:out = 10'b0010100011;        //489/3=163
			12'b000111101010:out = 10'b0010100011;        //490/3=163
			12'b000111101011:out = 10'b0010100011;        //491/3=163
			12'b000111101100:out = 10'b0010100100;        //492/3=164
			12'b000111101101:out = 10'b0010100100;        //493/3=164
			12'b000111101110:out = 10'b0010100100;        //494/3=164
			12'b000111101111:out = 10'b0010100101;        //495/3=165
			12'b000111110000:out = 10'b0010100101;        //496/3=165
			12'b000111110001:out = 10'b0010100101;        //497/3=165
			12'b000111110010:out = 10'b0010100110;        //498/3=166
			12'b000111110011:out = 10'b0010100110;        //499/3=166
			12'b000111110100:out = 10'b0010100110;        //500/3=166
			12'b000111110101:out = 10'b0010100111;        //501/3=167
			12'b000111110110:out = 10'b0010100111;        //502/3=167
			12'b000111110111:out = 10'b0010100111;        //503/3=167
			12'b000111111000:out = 10'b0010101000;        //504/3=168
			12'b000111111001:out = 10'b0010101000;        //505/3=168
			12'b000111111010:out = 10'b0010101000;        //506/3=168
			12'b000111111011:out = 10'b0010101001;        //507/3=169
			12'b000111111100:out = 10'b0010101001;        //508/3=169
			12'b000111111101:out = 10'b0010101001;        //509/3=169
			12'b000111111110:out = 10'b0010101010;        //510/3=170
			12'b000111111111:out = 10'b0010101010;        //511/3=170
			12'b001000000000:out = 10'b0010101010;        //512/3=170
			12'b001000000001:out = 10'b0010101011;        //513/3=171
			12'b001000000010:out = 10'b0010101011;        //514/3=171
			12'b001000000011:out = 10'b0010101011;        //515/3=171
			12'b001000000100:out = 10'b0010101100;        //516/3=172
			12'b001000000101:out = 10'b0010101100;        //517/3=172
			12'b001000000110:out = 10'b0010101100;        //518/3=172
			12'b001000000111:out = 10'b0010101101;        //519/3=173
			12'b001000001000:out = 10'b0010101101;        //520/3=173
			12'b001000001001:out = 10'b0010101101;        //521/3=173
			12'b001000001010:out = 10'b0010101110;        //522/3=174
			12'b001000001011:out = 10'b0010101110;        //523/3=174
			12'b001000001100:out = 10'b0010101110;        //524/3=174
			12'b001000001101:out = 10'b0010101111;        //525/3=175
			12'b001000001110:out = 10'b0010101111;        //526/3=175
			12'b001000001111:out = 10'b0010101111;        //527/3=175
			12'b001000010000:out = 10'b0010110000;        //528/3=176
			12'b001000010001:out = 10'b0010110000;        //529/3=176
			12'b001000010010:out = 10'b0010110000;        //530/3=176
			12'b001000010011:out = 10'b0010110001;        //531/3=177
			12'b001000010100:out = 10'b0010110001;        //532/3=177
			12'b001000010101:out = 10'b0010110001;        //533/3=177
			12'b001000010110:out = 10'b0010110010;        //534/3=178
			12'b001000010111:out = 10'b0010110010;        //535/3=178
			12'b001000011000:out = 10'b0010110010;        //536/3=178
			12'b001000011001:out = 10'b0010110011;        //537/3=179
			12'b001000011010:out = 10'b0010110011;        //538/3=179
			12'b001000011011:out = 10'b0010110011;        //539/3=179
			12'b001000011100:out = 10'b0010110100;        //540/3=180
			12'b001000011101:out = 10'b0010110100;        //541/3=180
			12'b001000011110:out = 10'b0010110100;        //542/3=180
			12'b001000011111:out = 10'b0010110101;        //543/3=181
			12'b001000100000:out = 10'b0010110101;        //544/3=181
			12'b001000100001:out = 10'b0010110101;        //545/3=181
			12'b001000100010:out = 10'b0010110110;        //546/3=182
			12'b001000100011:out = 10'b0010110110;        //547/3=182
			12'b001000100100:out = 10'b0010110110;        //548/3=182
			12'b001000100101:out = 10'b0010110111;        //549/3=183
			12'b001000100110:out = 10'b0010110111;        //550/3=183
			12'b001000100111:out = 10'b0010110111;        //551/3=183
			12'b001000101000:out = 10'b0010111000;        //552/3=184
			12'b001000101001:out = 10'b0010111000;        //553/3=184
			12'b001000101010:out = 10'b0010111000;        //554/3=184
			12'b001000101011:out = 10'b0010111001;        //555/3=185
			12'b001000101100:out = 10'b0010111001;        //556/3=185
			12'b001000101101:out = 10'b0010111001;        //557/3=185
			12'b001000101110:out = 10'b0010111010;        //558/3=186
			12'b001000101111:out = 10'b0010111010;        //559/3=186
			12'b001000110000:out = 10'b0010111010;        //560/3=186
			12'b001000110001:out = 10'b0010111011;        //561/3=187
			12'b001000110010:out = 10'b0010111011;        //562/3=187
			12'b001000110011:out = 10'b0010111011;        //563/3=187
			12'b001000110100:out = 10'b0010111100;        //564/3=188
			12'b001000110101:out = 10'b0010111100;        //565/3=188
			12'b001000110110:out = 10'b0010111100;        //566/3=188
			12'b001000110111:out = 10'b0010111101;        //567/3=189
			12'b001000111000:out = 10'b0010111101;        //568/3=189
			12'b001000111001:out = 10'b0010111101;        //569/3=189
			12'b001000111010:out = 10'b0010111110;        //570/3=190
			12'b001000111011:out = 10'b0010111110;        //571/3=190
			12'b001000111100:out = 10'b0010111110;        //572/3=190
			12'b001000111101:out = 10'b0010111111;        //573/3=191
			12'b001000111110:out = 10'b0010111111;        //574/3=191
			12'b001000111111:out = 10'b0010111111;        //575/3=191
			12'b001001000000:out = 10'b0011000000;        //576/3=192
			12'b001001000001:out = 10'b0011000000;        //577/3=192
			12'b001001000010:out = 10'b0011000000;        //578/3=192
			12'b001001000011:out = 10'b0011000001;        //579/3=193
			12'b001001000100:out = 10'b0011000001;        //580/3=193
			12'b001001000101:out = 10'b0011000001;        //581/3=193
			12'b001001000110:out = 10'b0011000010;        //582/3=194
			12'b001001000111:out = 10'b0011000010;        //583/3=194
			12'b001001001000:out = 10'b0011000010;        //584/3=194
			12'b001001001001:out = 10'b0011000011;        //585/3=195
			12'b001001001010:out = 10'b0011000011;        //586/3=195
			12'b001001001011:out = 10'b0011000011;        //587/3=195
			12'b001001001100:out = 10'b0011000100;        //588/3=196
			12'b001001001101:out = 10'b0011000100;        //589/3=196
			12'b001001001110:out = 10'b0011000100;        //590/3=196
			12'b001001001111:out = 10'b0011000101;        //591/3=197
			12'b001001010000:out = 10'b0011000101;        //592/3=197
			12'b001001010001:out = 10'b0011000101;        //593/3=197
			12'b001001010010:out = 10'b0011000110;        //594/3=198
			12'b001001010011:out = 10'b0011000110;        //595/3=198
			12'b001001010100:out = 10'b0011000110;        //596/3=198
			12'b001001010101:out = 10'b0011000111;        //597/3=199
			12'b001001010110:out = 10'b0011000111;        //598/3=199
			12'b001001010111:out = 10'b0011000111;        //599/3=199
			12'b001001011000:out = 10'b0011001000;        //600/3=200
			12'b001001011001:out = 10'b0011001000;        //601/3=200
			12'b001001011010:out = 10'b0011001000;        //602/3=200
			12'b001001011011:out = 10'b0011001001;        //603/3=201
			12'b001001011100:out = 10'b0011001001;        //604/3=201
			12'b001001011101:out = 10'b0011001001;        //605/3=201
			12'b001001011110:out = 10'b0011001010;        //606/3=202
			12'b001001011111:out = 10'b0011001010;        //607/3=202
			12'b001001100000:out = 10'b0011001010;        //608/3=202
			12'b001001100001:out = 10'b0011001011;        //609/3=203
			12'b001001100010:out = 10'b0011001011;        //610/3=203
			12'b001001100011:out = 10'b0011001011;        //611/3=203
			12'b001001100100:out = 10'b0011001100;        //612/3=204
			12'b001001100101:out = 10'b0011001100;        //613/3=204
			12'b001001100110:out = 10'b0011001100;        //614/3=204
			12'b001001100111:out = 10'b0011001101;        //615/3=205
			12'b001001101000:out = 10'b0011001101;        //616/3=205
			12'b001001101001:out = 10'b0011001101;        //617/3=205
			12'b001001101010:out = 10'b0011001110;        //618/3=206
			12'b001001101011:out = 10'b0011001110;        //619/3=206
			12'b001001101100:out = 10'b0011001110;        //620/3=206
			12'b001001101101:out = 10'b0011001111;        //621/3=207
			12'b001001101110:out = 10'b0011001111;        //622/3=207
			12'b001001101111:out = 10'b0011001111;        //623/3=207
			12'b001001110000:out = 10'b0011010000;        //624/3=208
			12'b001001110001:out = 10'b0011010000;        //625/3=208
			12'b001001110010:out = 10'b0011010000;        //626/3=208
			12'b001001110011:out = 10'b0011010001;        //627/3=209
			12'b001001110100:out = 10'b0011010001;        //628/3=209
			12'b001001110101:out = 10'b0011010001;        //629/3=209
			12'b001001110110:out = 10'b0011010010;        //630/3=210
			12'b001001110111:out = 10'b0011010010;        //631/3=210
			12'b001001111000:out = 10'b0011010010;        //632/3=210
			12'b001001111001:out = 10'b0011010011;        //633/3=211
			12'b001001111010:out = 10'b0011010011;        //634/3=211
			12'b001001111011:out = 10'b0011010011;        //635/3=211
			12'b001001111100:out = 10'b0011010100;        //636/3=212
			12'b001001111101:out = 10'b0011010100;        //637/3=212
			12'b001001111110:out = 10'b0011010100;        //638/3=212
			12'b001001111111:out = 10'b0011010101;        //639/3=213
			12'b001010000000:out = 10'b0011010101;        //640/3=213
			12'b001010000001:out = 10'b0011010101;        //641/3=213
			12'b001010000010:out = 10'b0011010110;        //642/3=214
			12'b001010000011:out = 10'b0011010110;        //643/3=214
			12'b001010000100:out = 10'b0011010110;        //644/3=214
			12'b001010000101:out = 10'b0011010111;        //645/3=215
			12'b001010000110:out = 10'b0011010111;        //646/3=215
			12'b001010000111:out = 10'b0011010111;        //647/3=215
			12'b001010001000:out = 10'b0011011000;        //648/3=216
			12'b001010001001:out = 10'b0011011000;        //649/3=216
			12'b001010001010:out = 10'b0011011000;        //650/3=216
			12'b001010001011:out = 10'b0011011001;        //651/3=217
			12'b001010001100:out = 10'b0011011001;        //652/3=217
			12'b001010001101:out = 10'b0011011001;        //653/3=217
			12'b001010001110:out = 10'b0011011010;        //654/3=218
			12'b001010001111:out = 10'b0011011010;        //655/3=218
			12'b001010010000:out = 10'b0011011010;        //656/3=218
			12'b001010010001:out = 10'b0011011011;        //657/3=219
			12'b001010010010:out = 10'b0011011011;        //658/3=219
			12'b001010010011:out = 10'b0011011011;        //659/3=219
			12'b001010010100:out = 10'b0011011100;        //660/3=220
			12'b001010010101:out = 10'b0011011100;        //661/3=220
			12'b001010010110:out = 10'b0011011100;        //662/3=220
			12'b001010010111:out = 10'b0011011101;        //663/3=221
			12'b001010011000:out = 10'b0011011101;        //664/3=221
			12'b001010011001:out = 10'b0011011101;        //665/3=221
			12'b001010011010:out = 10'b0011011110;        //666/3=222
			12'b001010011011:out = 10'b0011011110;        //667/3=222
			12'b001010011100:out = 10'b0011011110;        //668/3=222
			12'b001010011101:out = 10'b0011011111;        //669/3=223
			12'b001010011110:out = 10'b0011011111;        //670/3=223
			12'b001010011111:out = 10'b0011011111;        //671/3=223
			12'b001010100000:out = 10'b0011100000;        //672/3=224
			12'b001010100001:out = 10'b0011100000;        //673/3=224
			12'b001010100010:out = 10'b0011100000;        //674/3=224
			12'b001010100011:out = 10'b0011100001;        //675/3=225
			12'b001010100100:out = 10'b0011100001;        //676/3=225
			12'b001010100101:out = 10'b0011100001;        //677/3=225
			12'b001010100110:out = 10'b0011100010;        //678/3=226
			12'b001010100111:out = 10'b0011100010;        //679/3=226
			12'b001010101000:out = 10'b0011100010;        //680/3=226
			12'b001010101001:out = 10'b0011100011;        //681/3=227
			12'b001010101010:out = 10'b0011100011;        //682/3=227
			12'b001010101011:out = 10'b0011100011;        //683/3=227
			12'b001010101100:out = 10'b0011100100;        //684/3=228
			12'b001010101101:out = 10'b0011100100;        //685/3=228
			12'b001010101110:out = 10'b0011100100;        //686/3=228
			12'b001010101111:out = 10'b0011100101;        //687/3=229
			12'b001010110000:out = 10'b0011100101;        //688/3=229
			12'b001010110001:out = 10'b0011100101;        //689/3=229
			12'b001010110010:out = 10'b0011100110;        //690/3=230
			12'b001010110011:out = 10'b0011100110;        //691/3=230
			12'b001010110100:out = 10'b0011100110;        //692/3=230
			12'b001010110101:out = 10'b0011100111;        //693/3=231
			12'b001010110110:out = 10'b0011100111;        //694/3=231
			12'b001010110111:out = 10'b0011100111;        //695/3=231
			12'b001010111000:out = 10'b0011101000;        //696/3=232
			12'b001010111001:out = 10'b0011101000;        //697/3=232
			12'b001010111010:out = 10'b0011101000;        //698/3=232
			12'b001010111011:out = 10'b0011101001;        //699/3=233
			12'b001010111100:out = 10'b0011101001;        //700/3=233
			12'b001010111101:out = 10'b0011101001;        //701/3=233
			12'b001010111110:out = 10'b0011101010;        //702/3=234
			12'b001010111111:out = 10'b0011101010;        //703/3=234
			12'b001011000000:out = 10'b0011101010;        //704/3=234
			12'b001011000001:out = 10'b0011101011;        //705/3=235
			12'b001011000010:out = 10'b0011101011;        //706/3=235
			12'b001011000011:out = 10'b0011101011;        //707/3=235
			12'b001011000100:out = 10'b0011101100;        //708/3=236
			12'b001011000101:out = 10'b0011101100;        //709/3=236
			12'b001011000110:out = 10'b0011101100;        //710/3=236
			12'b001011000111:out = 10'b0011101101;        //711/3=237
			12'b001011001000:out = 10'b0011101101;        //712/3=237
			12'b001011001001:out = 10'b0011101101;        //713/3=237
			12'b001011001010:out = 10'b0011101110;        //714/3=238
			12'b001011001011:out = 10'b0011101110;        //715/3=238
			12'b001011001100:out = 10'b0011101110;        //716/3=238
			12'b001011001101:out = 10'b0011101111;        //717/3=239
			12'b001011001110:out = 10'b0011101111;        //718/3=239
			12'b001011001111:out = 10'b0011101111;        //719/3=239
			12'b001011010000:out = 10'b0011110000;        //720/3=240
			12'b001011010001:out = 10'b0011110000;        //721/3=240
			12'b001011010010:out = 10'b0011110000;        //722/3=240
			12'b001011010011:out = 10'b0011110001;        //723/3=241
			12'b001011010100:out = 10'b0011110001;        //724/3=241
			12'b001011010101:out = 10'b0011110001;        //725/3=241
			12'b001011010110:out = 10'b0011110010;        //726/3=242
			12'b001011010111:out = 10'b0011110010;        //727/3=242
			12'b001011011000:out = 10'b0011110010;        //728/3=242
			12'b001011011001:out = 10'b0011110011;        //729/3=243
			12'b001011011010:out = 10'b0011110011;        //730/3=243
			12'b001011011011:out = 10'b0011110011;        //731/3=243
			12'b001011011100:out = 10'b0011110100;        //732/3=244
			12'b001011011101:out = 10'b0011110100;        //733/3=244
			12'b001011011110:out = 10'b0011110100;        //734/3=244
			12'b001011011111:out = 10'b0011110101;        //735/3=245
			12'b001011100000:out = 10'b0011110101;        //736/3=245
			12'b001011100001:out = 10'b0011110101;        //737/3=245
			12'b001011100010:out = 10'b0011110110;        //738/3=246
			12'b001011100011:out = 10'b0011110110;        //739/3=246
			12'b001011100100:out = 10'b0011110110;        //740/3=246
			12'b001011100101:out = 10'b0011110111;        //741/3=247
			12'b001011100110:out = 10'b0011110111;        //742/3=247
			12'b001011100111:out = 10'b0011110111;        //743/3=247
			12'b001011101000:out = 10'b0011111000;        //744/3=248
			12'b001011101001:out = 10'b0011111000;        //745/3=248
			12'b001011101010:out = 10'b0011111000;        //746/3=248
			12'b001011101011:out = 10'b0011111001;        //747/3=249
			12'b001011101100:out = 10'b0011111001;        //748/3=249
			12'b001011101101:out = 10'b0011111001;        //749/3=249
			12'b001011101110:out = 10'b0011111010;        //750/3=250
			12'b001011101111:out = 10'b0011111010;        //751/3=250
			12'b001011110000:out = 10'b0011111010;        //752/3=250
			12'b001011110001:out = 10'b0011111011;        //753/3=251
			12'b001011110010:out = 10'b0011111011;        //754/3=251
			12'b001011110011:out = 10'b0011111011;        //755/3=251
			12'b001011110100:out = 10'b0011111100;        //756/3=252
			12'b001011110101:out = 10'b0011111100;        //757/3=252
			12'b001011110110:out = 10'b0011111100;        //758/3=252
			12'b001011110111:out = 10'b0011111101;        //759/3=253
			12'b001011111000:out = 10'b0011111101;        //760/3=253
			12'b001011111001:out = 10'b0011111101;        //761/3=253
			12'b001011111010:out = 10'b0011111110;        //762/3=254
			12'b001011111011:out = 10'b0011111110;        //763/3=254
			12'b001011111100:out = 10'b0011111110;        //764/3=254
			12'b001011111101:out = 10'b0011111111;        //765/3=255
			12'b001011111110:out = 10'b0011111111;        //766/3=255
			12'b001011111111:out = 10'b0011111111;        //767/3=255
			12'b001100000000:out = 10'b0100000000;        //768/3=256
			12'b001100000001:out = 10'b0100000000;        //769/3=256
			12'b001100000010:out = 10'b0100000000;        //770/3=256
			12'b001100000011:out = 10'b0100000001;        //771/3=257
			12'b001100000100:out = 10'b0100000001;        //772/3=257
			12'b001100000101:out = 10'b0100000001;        //773/3=257
			12'b001100000110:out = 10'b0100000010;        //774/3=258
			12'b001100000111:out = 10'b0100000010;        //775/3=258
			12'b001100001000:out = 10'b0100000010;        //776/3=258
			12'b001100001001:out = 10'b0100000011;        //777/3=259
			12'b001100001010:out = 10'b0100000011;        //778/3=259
			12'b001100001011:out = 10'b0100000011;        //779/3=259
			12'b001100001100:out = 10'b0100000100;        //780/3=260
			12'b001100001101:out = 10'b0100000100;        //781/3=260
			12'b001100001110:out = 10'b0100000100;        //782/3=260
			12'b001100001111:out = 10'b0100000101;        //783/3=261
			12'b001100010000:out = 10'b0100000101;        //784/3=261
			12'b001100010001:out = 10'b0100000101;        //785/3=261
			12'b001100010010:out = 10'b0100000110;        //786/3=262
			12'b001100010011:out = 10'b0100000110;        //787/3=262
			12'b001100010100:out = 10'b0100000110;        //788/3=262
			12'b001100010101:out = 10'b0100000111;        //789/3=263
			12'b001100010110:out = 10'b0100000111;        //790/3=263
			12'b001100010111:out = 10'b0100000111;        //791/3=263
			12'b001100011000:out = 10'b0100001000;        //792/3=264
			12'b001100011001:out = 10'b0100001000;        //793/3=264
			12'b001100011010:out = 10'b0100001000;        //794/3=264
			12'b001100011011:out = 10'b0100001001;        //795/3=265
			12'b001100011100:out = 10'b0100001001;        //796/3=265
			12'b001100011101:out = 10'b0100001001;        //797/3=265
			12'b001100011110:out = 10'b0100001010;        //798/3=266
			12'b001100011111:out = 10'b0100001010;        //799/3=266
			12'b001100100000:out = 10'b0100001010;        //800/3=266
			12'b001100100001:out = 10'b0100001011;        //801/3=267
			12'b001100100010:out = 10'b0100001011;        //802/3=267
			12'b001100100011:out = 10'b0100001011;        //803/3=267
			12'b001100100100:out = 10'b0100001100;        //804/3=268
			12'b001100100101:out = 10'b0100001100;        //805/3=268
			12'b001100100110:out = 10'b0100001100;        //806/3=268
			12'b001100100111:out = 10'b0100001101;        //807/3=269
			12'b001100101000:out = 10'b0100001101;        //808/3=269
			12'b001100101001:out = 10'b0100001101;        //809/3=269
			12'b001100101010:out = 10'b0100001110;        //810/3=270
			12'b001100101011:out = 10'b0100001110;        //811/3=270
			12'b001100101100:out = 10'b0100001110;        //812/3=270
			12'b001100101101:out = 10'b0100001111;        //813/3=271
			12'b001100101110:out = 10'b0100001111;        //814/3=271
			12'b001100101111:out = 10'b0100001111;        //815/3=271
			12'b001100110000:out = 10'b0100010000;        //816/3=272
			12'b001100110001:out = 10'b0100010000;        //817/3=272
			12'b001100110010:out = 10'b0100010000;        //818/3=272
			12'b001100110011:out = 10'b0100010001;        //819/3=273
			12'b001100110100:out = 10'b0100010001;        //820/3=273
			12'b001100110101:out = 10'b0100010001;        //821/3=273
			12'b001100110110:out = 10'b0100010010;        //822/3=274
			12'b001100110111:out = 10'b0100010010;        //823/3=274
			12'b001100111000:out = 10'b0100010010;        //824/3=274
			12'b001100111001:out = 10'b0100010011;        //825/3=275
			12'b001100111010:out = 10'b0100010011;        //826/3=275
			12'b001100111011:out = 10'b0100010011;        //827/3=275
			12'b001100111100:out = 10'b0100010100;        //828/3=276
			12'b001100111101:out = 10'b0100010100;        //829/3=276
			12'b001100111110:out = 10'b0100010100;        //830/3=276
			12'b001100111111:out = 10'b0100010101;        //831/3=277
			12'b001101000000:out = 10'b0100010101;        //832/3=277
			12'b001101000001:out = 10'b0100010101;        //833/3=277
			12'b001101000010:out = 10'b0100010110;        //834/3=278
			12'b001101000011:out = 10'b0100010110;        //835/3=278
			12'b001101000100:out = 10'b0100010110;        //836/3=278
			12'b001101000101:out = 10'b0100010111;        //837/3=279
			12'b001101000110:out = 10'b0100010111;        //838/3=279
			12'b001101000111:out = 10'b0100010111;        //839/3=279
			12'b001101001000:out = 10'b0100011000;        //840/3=280
			12'b001101001001:out = 10'b0100011000;        //841/3=280
			12'b001101001010:out = 10'b0100011000;        //842/3=280
			12'b001101001011:out = 10'b0100011001;        //843/3=281
			12'b001101001100:out = 10'b0100011001;        //844/3=281
			12'b001101001101:out = 10'b0100011001;        //845/3=281
			12'b001101001110:out = 10'b0100011010;        //846/3=282
			12'b001101001111:out = 10'b0100011010;        //847/3=282
			12'b001101010000:out = 10'b0100011010;        //848/3=282
			12'b001101010001:out = 10'b0100011011;        //849/3=283
			12'b001101010010:out = 10'b0100011011;        //850/3=283
			12'b001101010011:out = 10'b0100011011;        //851/3=283
			12'b001101010100:out = 10'b0100011100;        //852/3=284
			12'b001101010101:out = 10'b0100011100;        //853/3=284
			12'b001101010110:out = 10'b0100011100;        //854/3=284
			12'b001101010111:out = 10'b0100011101;        //855/3=285
			12'b001101011000:out = 10'b0100011101;        //856/3=285
			12'b001101011001:out = 10'b0100011101;        //857/3=285
			12'b001101011010:out = 10'b0100011110;        //858/3=286
			12'b001101011011:out = 10'b0100011110;        //859/3=286
			12'b001101011100:out = 10'b0100011110;        //860/3=286
			12'b001101011101:out = 10'b0100011111;        //861/3=287 
			12'b001101011110:out = 10'b0100011111;        //862/3=287
			12'b001101011111:out = 10'b0100011111;        //863/3=287
			12'b001101100000:out = 10'b0100100000;        //864/3=288
			12'b001101100001:out = 10'b0100100000;        //865/3=288
			12'b001101100010:out = 10'b0100100000;        //866/3=288
			12'b001101100011:out = 10'b0100100001;        //867/3=289
			12'b001101100100:out = 10'b0100100001;        //868/3=289
			12'b001101100101:out = 10'b0100100001;        //869/3=289
			12'b001101100110:out = 10'b0100100010;        //870/3=290
			12'b001101100111:out = 10'b0100100010;        //871/3=290
			12'b001101101000:out = 10'b0100100010;        //872/3=290
			12'b001101101001:out = 10'b0100100011;        //873/3=291
			12'b001101101010:out = 10'b0100100011;        //874/3=291
			12'b001101101011:out = 10'b0100100011;        //875/3=291
			12'b001101101100:out = 10'b0100100100;        //876/3=292
			12'b001101101101:out = 10'b0100100100;        //877/3=292
			12'b001101101110:out = 10'b0100100100;        //878/3=292
			12'b001101101111:out = 10'b0100100101;        //879/3=293
			12'b001101110000:out = 10'b0100100101;        //880/3=293
			12'b001101110001:out = 10'b0100100101;        //881/3=293
			12'b001101110010:out = 10'b0100100110;        //882/3=294
			12'b001101110011:out = 10'b0100100110;        //883/3=294
			12'b001101110100:out = 10'b0100100110;        //884/3=294
			12'b001101110101:out = 10'b0100100111;        //885/3=295
			12'b001101110110:out = 10'b0100100111;        //886/3=295
			12'b001101110111:out = 10'b0100100111;        //887/3=295
			12'b001101111000:out = 10'b0100101000;        //888/3=296
			12'b001101111001:out = 10'b0100101000;        //889/3=296
			12'b001101111010:out = 10'b0100101000;        //890/3=296
			12'b001101111011:out = 10'b0100101001;        //891/3=297
			12'b001101111100:out = 10'b0100101001;        //892/3=297
			12'b001101111101:out = 10'b0100101001;        //893/3=297
			12'b001101111110:out = 10'b0100101010;        //894/3=298
			12'b001101111111:out = 10'b0100101010;        //895/3=298
			12'b001110000000:out = 10'b0100101010;        //896/3=298
			12'b001110000001:out = 10'b0100101011;        //897/3=299
			12'b001110000010:out = 10'b0100101011;        //898/3=299
			12'b001110000011:out = 10'b0100101011;        //899/3=299
			12'b001110000100:out = 10'b0100101100;        //900/3=300
			12'b001110000101:out = 10'b0100101100;        //901/3=300
			12'b001110000110:out = 10'b0100101100;        //902/3=300
			12'b001110000111:out = 10'b0100101101;        //903/3=301
			12'b001110001000:out = 10'b0100101101;        //904/3=301
			12'b001110001001:out = 10'b0100101101;        //905/3=301
			12'b001110001010:out = 10'b0100101110;        //906/3=302
			12'b001110001011:out = 10'b0100101110;        //907/3=302
			12'b001110001100:out = 10'b0100101110;        //908/3=302
			12'b001110001101:out = 10'b0100101111;        //909/3=303
			12'b001110001110:out = 10'b0100101111;        //910/3=303
			12'b001110001111:out = 10'b0100101111;        //911/3=303
			12'b001110010000:out = 10'b0100110000;        //912/3=304
			12'b001110010001:out = 10'b0100110000;        //913/3=304
			12'b001110010010:out = 10'b0100110000;        //914/3=304
			12'b001110010011:out = 10'b0100110001;        //915/3=305
			12'b001110010100:out = 10'b0100110001;        //916/3=305
			12'b001110010101:out = 10'b0100110001;        //917/3=305
			12'b001110010110:out = 10'b0100110010;        //918/3=306
			12'b001110010111:out = 10'b0100110010;        //919/3=306
			12'b001110011000:out = 10'b0100110010;        //920/3=306
			12'b001110011001:out = 10'b0100110011;        //921/3=307
			12'b001110011010:out = 10'b0100110011;        //922/3=307
			12'b001110011011:out = 10'b0100110011;        //923/3=307
			12'b001110011100:out = 10'b0100110100;        //924/3=308
			12'b001110011101:out = 10'b0100110100;        //925/3=308
			12'b001110011110:out = 10'b0100110100;        //926/3=308
			12'b001110011111:out = 10'b0100110101;        //927/3=309
			12'b001110100000:out = 10'b0100110101;        //928/3=309
			12'b001110100001:out = 10'b0100110101;        //929/3=309
			12'b001110100010:out = 10'b0100110110;        //930/3=310
			12'b001110100011:out = 10'b0100110110;        //931/3=310
			12'b001110100100:out = 10'b0100110110;        //932/3=310
			12'b001110100101:out = 10'b0100110111;        //933/3=311
			12'b001110100110:out = 10'b0100110111;        //934/3=311
			12'b001110100111:out = 10'b0100110111;        //935/3=311
			12'b001110101000:out = 10'b0100111000;        //936/3=312
			12'b001110101001:out = 10'b0100111000;        //937/3=312
			12'b001110101010:out = 10'b0100111000;        //938/3=312
			12'b001110101011:out = 10'b0100111001;        //939/3=313
			12'b001110101100:out = 10'b0100111001;        //940/3=313
			12'b001110101101:out = 10'b0100111001;        //941/3=313
			12'b001110101110:out = 10'b0100111010;        //942/3=314
			12'b001110101111:out = 10'b0100111010;        //943/3=314
			12'b001110110000:out = 10'b0100111010;        //944/3=314
			12'b001110110001:out = 10'b0100111011;        //945/3=315
			12'b001110110010:out = 10'b0100111011;        //946/3=315
			12'b001110110011:out = 10'b0100111011;        //947/3=315
			12'b001110110100:out = 10'b0100111100;        //948/3=316
			12'b001110110101:out = 10'b0100111100;        //949/3=316
			12'b001110110110:out = 10'b0100111100;        //950/3=316
			12'b001110110111:out = 10'b0100111101;        //951/3=317
			12'b001110111000:out = 10'b0100111101;        //952/3=317
			12'b001110111001:out = 10'b0100111101;        //953/3=317
			12'b001110111010:out = 10'b0100111110;        //954/3=318
			12'b001110111011:out = 10'b0100111110;        //955/3=318
			12'b001110111100:out = 10'b0100111110;        //956/3=318
			12'b001110111101:out = 10'b0100111111;        //957/3=319
			12'b001110111110:out = 10'b0100111111;        //958/3=319
			12'b001110111111:out = 10'b0100111111;        //959/3=319
			12'b001111000000:out = 10'b0101000000;        //960/3=320
			12'b001111000001:out = 10'b0101000000;        //961/3=320
			12'b001111000010:out = 10'b0101000000;        //962/3=320
			12'b001111000011:out = 10'b0101000001;        //963/3=321
			12'b001111000100:out = 10'b0101000001;        //964/3=321
			12'b001111000101:out = 10'b0101000001;        //965/3=321
			12'b001111000110:out = 10'b0101000010;        //966/3=322
			12'b001111000111:out = 10'b0101000010;        //967/3=322
			12'b001111001000:out = 10'b0101000010;        //968/3=322
			12'b001111001001:out = 10'b0101000011;        //969/3=323
			12'b001111001010:out = 10'b0101000011;        //970/3=323
			12'b001111001011:out = 10'b0101000011;        //971/3=323
			12'b001111001100:out = 10'b0101000100;        //972/3=324
			12'b001111001101:out = 10'b0101000100;        //973/3=324
			12'b001111001110:out = 10'b0101000100;        //974/3=324
			12'b001111001111:out = 10'b0101000101;        //975/3=325
			12'b001111010000:out = 10'b0101000101;        //976/3=325
			12'b001111010001:out = 10'b0101000101;        //977/3=325
			12'b001111010010:out = 10'b0101000110;        //978/3=326
			12'b001111010011:out = 10'b0101000110;        //979/3=326
			12'b001111010100:out = 10'b0101000110;        //980/3=326
			12'b001111010101:out = 10'b0101000111;        //981/3=327
			12'b001111010110:out = 10'b0101000111;        //982/3=327
			12'b001111010111:out = 10'b0101000111;        //983/3=327
			12'b001111011000:out = 10'b0101001000;        //984/3=328
			12'b001111011001:out = 10'b0101001000;        //985/3=328
			12'b001111011010:out = 10'b0101001000;        //986/3=328
			12'b001111011011:out = 10'b0101001001;        //987/3=329
			12'b001111011100:out = 10'b0101001001;        //988/3=329
			12'b001111011101:out = 10'b0101001001;        //989/3=329
			12'b001111011110:out = 10'b0101001010;        //990/3=330
			12'b001111011111:out = 10'b0101001010;        //991/3=330
			12'b001111100000:out = 10'b0101001010;        //992/3=330
			12'b001111100001:out = 10'b0101001011;        //993/3=331
			12'b001111100010:out = 10'b0101001011;        //994/3=331
			12'b001111100011:out = 10'b0101001011;        //995/3=331
			12'b001111100100:out = 10'b0101001100;        //996/3=332
			12'b001111100101:out = 10'b0101001100;        //997/3=332
			12'b001111100110:out = 10'b0101001100;        //998/3=332
			12'b001111100111:out = 10'b0101001101;        //999/3=333
			12'b001111101000:out = 10'b0101001101;        //1000/3=333
			12'b001111101001:out = 10'b0101001101;        //1001/3=333
			12'b001111101010:out = 10'b0101001110;        //1002/3=334
			12'b001111101011:out = 10'b0101001110;        //1003/3=334
			12'b001111101100:out = 10'b0101001110;        //1004/3=334
			12'b001111101101:out = 10'b0101001111;        //1005/3=335
			12'b001111101110:out = 10'b0101001111;        //1006/3=335
			12'b001111101111:out = 10'b0101001111;        //1007/3=335
			12'b001111110000:out = 10'b0101010000;        //1008/3=336
			12'b001111110001:out = 10'b0101010000;        //1009/3=336
			12'b001111110010:out = 10'b0101010000;        //1010/3=336
			12'b001111110011:out = 10'b0101010001;        //1011/3=337
			12'b001111110100:out = 10'b0101010001;        //1012/3=337
			12'b001111110101:out = 10'b0101010001;        //1013/3=337
			12'b001111110110:out = 10'b0101010010;        //1014/3=338
			12'b001111110111:out = 10'b0101010010;        //1015/3=338
			12'b001111111000:out = 10'b0101010010;        //1016/3=338
			12'b001111111001:out = 10'b0101010011;        //1017/3=339
			12'b001111111010:out = 10'b0101010011;        //1018/3=339
			12'b001111111011:out = 10'b0101010011;        //1019/3=339
			12'b001111111100:out = 10'b0101010100;        //1020/3=340
			12'b001111111101:out = 10'b0101010100;        //1021/3=340
			12'b001111111110:out = 10'b0101010100;        //1022/3=340
			12'b001111111111:out = 10'b0101010101;        //1023/3=341
			12'b010000000000:out = 10'b0101010101;        //1024/3=341
			12'b010000000001:out = 10'b0101010101;        //1025/3=341
			12'b010000000010:out = 10'b0101010110;        //1026/3=342
			12'b010000000011:out = 10'b0101010110;        //1027/3=342
			12'b010000000100:out = 10'b0101010110;        //1028/3=342
			12'b010000000101:out = 10'b0101010111;        //1029/3=343
			12'b010000000110:out = 10'b0101010111;        //1030/3=343
			12'b010000000111:out = 10'b0101010111;        //1031/3=343
			12'b010000001000:out = 10'b0101011000;        //1032/3=344
			12'b010000001001:out = 10'b0101011000;        //1033/3=344
			12'b010000001010:out = 10'b0101011000;        //1034/3=344
			12'b010000001011:out = 10'b0101011001;        //1035/3=345
			12'b010000001100:out = 10'b0101011001;        //1036/3=345
			12'b010000001101:out = 10'b0101011001;        //1037/3=345
			12'b010000001110:out = 10'b0101011010;        //1038/3=346
			12'b010000001111:out = 10'b0101011010;        //1039/3=346
			12'b010000010000:out = 10'b0101011010;        //1040/3=346
			12'b010000010001:out = 10'b0101011011;        //1041/3=347
			12'b010000010010:out = 10'b0101011011;        //1042/3=347
			12'b010000010011:out = 10'b0101011011;        //1043/3=347
			12'b010000010100:out = 10'b0101011100;        //1044/3=348
			12'b010000010101:out = 10'b0101011100;        //1045/3=348
			12'b010000010110:out = 10'b0101011100;        //1046/3=348
			12'b010000010111:out = 10'b0101011101;        //1047/3=349
			12'b010000011000:out = 10'b0101011101;        //1048/3=349
			12'b010000011001:out = 10'b0101011101;        //1049/3=349
			12'b010000011010:out = 10'b0101011110;        //1050/3=350
			12'b010000011011:out = 10'b0101011110;        //1051/3=350
			12'b010000011100:out = 10'b0101011110;        //1052/3=350
			12'b010000011101:out = 10'b0101011111;        //1053/3=351
			12'b010000011110:out = 10'b0101011111;        //1054/3=351
			12'b010000011111:out = 10'b0101011111;        //1055/3=351
			12'b010000100000:out = 10'b0101100000;        //1056/3=352
			12'b010000100001:out = 10'b0101100000;        //1057/3=352
			12'b010000100010:out = 10'b0101100000;        //1058/3=352
			12'b010000100011:out = 10'b0101100001;        //1059/3=353
			12'b010000100100:out = 10'b0101100001;        //1060/3=353
			12'b010000100101:out = 10'b0101100001;        //1061/3=353
			12'b010000100110:out = 10'b0101100010;        //1062/3=354
			12'b010000100111:out = 10'b0101100010;        //1063/3=354
			12'b010000101000:out = 10'b0101100010;        //1064/3=354
			12'b010000101001:out = 10'b0101100011;        //1065/3=355
			12'b010000101010:out = 10'b0101100011;        //1066/3=355
			12'b010000101011:out = 10'b0101100011;        //1067/3=355
			12'b010000101100:out = 10'b0101100100;        //1068/3=356
			12'b010000101101:out = 10'b0101100100;        //1069/3=356
			12'b010000101110:out = 10'b0101100100;        //1070/3=356
			12'b010000101111:out = 10'b0101100101;        //1071/3=357
			12'b010000110000:out = 10'b0101100101;        //1072/3=357
			12'b010000110001:out = 10'b0101100101;        //1073/3=357
			12'b010000110010:out = 10'b0101100110;        //1074/3=358
			12'b010000110011:out = 10'b0101100110;        //1075/3=358
			12'b010000110100:out = 10'b0101100110;        //1076/3=358
			12'b010000110101:out = 10'b0101100111;        //1077/3=359
			12'b010000110110:out = 10'b0101100111;        //1078/3=359
			12'b010000110111:out = 10'b0101100111;        //1079/3=359
			12'b010000111000:out = 10'b0101101000;        //1080/3=360
			12'b010000111001:out = 10'b0101101000;        //1081/3=360
			12'b010000111010:out = 10'b0101101000;        //1082/3=360
			12'b010000111011:out = 10'b0101101001;        //1083/3=361
			12'b010000111100:out = 10'b0101101001;        //1084/3=361
			12'b010000111101:out = 10'b0101101001;        //1085/3=361
			12'b010000111110:out = 10'b0101101010;        //1086/3=362
			12'b010000111111:out = 10'b0101101010;        //1087/3=362
			12'b010001000000:out = 10'b0101101010;        //1088/3=362
			12'b010001000001:out = 10'b0101101011;        //1089/3=363
			12'b010001000010:out = 10'b0101101011;        //1090/3=363
			12'b010001000011:out = 10'b0101101011;        //1091/3=363
			12'b010001000100:out = 10'b0101101100;        //1092/3=364
			12'b010001000101:out = 10'b0101101100;        //1093/3=364
			12'b010001000110:out = 10'b0101101100;        //1094/3=364
			12'b010001000111:out = 10'b0101101101;        //1095/3=365
			12'b010001001000:out = 10'b0101101101;        //1096/3=365
			12'b010001001001:out = 10'b0101101101;        //1097/3=365
			12'b010001001010:out = 10'b0101101110;        //1098/3=366
			12'b010001001011:out = 10'b0101101110;        //1099/3=366
			12'b010001001100:out = 10'b0101101110;        //1100/3=366
			12'b010001001101:out = 10'b0101101111;        //1101/3=367
			12'b010001001110:out = 10'b0101101111;        //1102/3=367
			12'b010001001111:out = 10'b0101101111;        //1103/3=367
			12'b010001010000:out = 10'b0101110000;        //1104/3=368
			12'b010001010001:out = 10'b0101110000;        //1105/3=368
			12'b010001010010:out = 10'b0101110000;        //1106/3=368
			12'b010001010011:out = 10'b0101110001;        //1107/3=369
			12'b010001010100:out = 10'b0101110001;        //1108/3=369
			12'b010001010101:out = 10'b0101110001;        //1109/3=369
			12'b010001010110:out = 10'b0101110010;        //1110/3=370
			12'b010001010111:out = 10'b0101110010;        //1111/3=370
			12'b010001011000:out = 10'b0101110010;        //1112/3=370
			12'b010001011001:out = 10'b0101110011;        //1113/3=371
			12'b010001011010:out = 10'b0101110011;        //1114/3=371
			12'b010001011011:out = 10'b0101110011;        //1115/3=371
			12'b010001011100:out = 10'b0101110100;        //1116/3=372
			12'b010001011101:out = 10'b0101110100;        //1117/3=372
			12'b010001011110:out = 10'b0101110100;        //1118/3=372
			12'b010001100000:out = 10'b0101110101;        //1120/3=373
			12'b010001100001:out = 10'b0101110101;        //1121/3=373
			12'b010001100010:out = 10'b0101110110;        //1122/3=374
			12'b010001100100:out = 10'b0101110110;        //1124/3=374
			12'b010001100101:out = 10'b0101110111;        //1125/3=375
			default:out = 10'bx;

		endcase
endmodule


module div_3(
	input [6:0]in,
	output reg[4:0]out
);
	always@(in)
		case(in)
			7'b0000000:out = 5'b00000;        //0/3=0
			7'b0000001:out = 5'b00000;        //1/3=0
			7'b0000010:out = 5'b00000;        //2/3=0
			7'b0000011:out = 5'b00001;        //3/3=1
			7'b0000100:out = 5'b00001;        //4/3=1
			7'b0000101:out = 5'b00001;        //5/3=1
			7'b0000110:out = 5'b00010;        //6/3=2
			7'b0000111:out = 5'b00010;        //7/3=2
			7'b0001000:out = 5'b00010;        //8/3=2
			7'b0001001:out = 5'b00011;        //9/3=3
			7'b0001010:out = 5'b00011;        //10/3=3
			7'b0001011:out = 5'b00011;        //11/3=3
			7'b0001100:out = 5'b00100;        //12/3=4
			7'b0001101:out = 5'b00100;        //13/3=4
			7'b0001110:out = 5'b00100;        //14/3=4
			7'b0001111:out = 5'b00101;        //15/3=5
			7'b0010000:out = 5'b00101;        //16/3=5
			7'b0010001:out = 5'b00101;        //17/3=5
			7'b0010010:out = 5'b00110;        //18/3=6
			7'b0010011:out = 5'b00110;        //19/3=6
			7'b0010100:out = 5'b00110;        //20/3=6
			7'b0010101:out = 5'b00111;        //21/3=7
			7'b0010110:out = 5'b00111;        //22/3=7
			7'b0010111:out = 5'b00111;        //23/3=7
			7'b0011000:out = 5'b01000;        //24/3=8
			7'b0011001:out = 5'b01000;        //25/3=8
			7'b0011010:out = 5'b01000;        //26/3=8
			7'b0011011:out = 5'b01001;        //27/3=9
			7'b0011100:out = 5'b01001;        //28/3=9
			7'b0011101:out = 5'b01001;        //29/3=9
			7'b0011110:out = 5'b01010;        //30/3=10
			7'b0011111:out = 5'b01010;        //31/3=10
			7'b0100000:out = 5'b01010;        //32/3=10
			7'b0100001:out = 5'b01011;        //33/3=11
			7'b0100010:out = 5'b01011;        //34/3=11
			7'b0100011:out = 5'b01011;        //35/3=11
			7'b0100100:out = 5'b01100;        //36/3=12
			7'b0100101:out = 5'b01100;        //37/3=12
			7'b0100110:out = 5'b01100;        //38/3=12
			7'b0100111:out = 5'b01101;        //39/3=13
			7'b0101000:out = 5'b01101;        //40/3=13
			7'b0101001:out = 5'b01101;        //41/3=13
			7'b0101010:out = 5'b01110;        //42/3=14
			7'b0101011:out = 5'b01110;        //43/3=14
			7'b0101100:out = 5'b01110;        //44/3=14
			7'b0101101:out = 5'b01111;        //45/3=15
			
			7'b1101000:out = 5'b11000;        //-24/3=-8
			7'b1101001:out = 5'b11001;        //-23/3=-7
			7'b1101010:out = 5'b11001;        //-22/3=-7
			7'b1101011:out = 5'b11001;        //-21/3=-7
			7'b1101100:out = 5'b11010;        //-20/3=-6
			7'b1101101:out = 5'b11010;        //-19/3=-6
			7'b1101110:out = 5'b11010;        //-18/3=-6
			7'b1101111:out = 5'b11011;        //-17/3=-5
			7'b1110000:out = 5'b11011;        //-16/3=-5
			7'b1110001:out = 5'b11011;        //-15/3=-5
			7'b1110010:out = 5'b11100;        //-14/3=-4
			7'b1110011:out = 5'b11100;        //-13/3=-4
			7'b1110100:out = 5'b11100;        //-12/3=-4
			7'b1110101:out = 5'b11101;        //-11/3=-3
			7'b1110110:out = 5'b11101;        //-10/3=-3
			7'b1110111:out = 5'b11101;        //-9/3=-3
			7'b1111000:out = 5'b11110;        //-8/3=-2
			7'b1111001:out = 5'b11110;        //-7/3=-2
			7'b1111010:out = 5'b11110;        //-6/3=-2
			7'b1111011:out = 5'b11111;        //-5/3=-1
			7'b1111100:out = 5'b11111;        //-4/3=-1
			7'b1111101:out = 5'b11111;        //-3/3=-1
			7'b1111110:out = 5'b00000;        //-2/3=0
			7'b1111111:out = 5'b00000;        //-1/3=0
			
			default   :out = 5'bx;
		endcase
endmodule


module CC(
	in_n0,
	in_n1, 
	in_n2, 
	in_n3, 
    in_n4, 
	in_n5, 
	opt,
    equ,
	out_n
);
input wire [3:0]in_n0;
input wire [3:0]in_n1;
input wire [3:0]in_n2;
input wire [3:0]in_n3;
input wire [3:0]in_n4;
input wire [3:0]in_n5;
input wire [2:0] opt;
input wire equ;
output wire [9:0] out_n;
//==================================================================
// reg & wire
//==================================================================
wire [3:0]node00,node01,node02,node03,node04,node05,	
	node10,node11,node12,node13,node14,node15,
	node21,node22,node23,node24,
	node32,node33;
	
wire [3:0]sorted0,sorted1,sorted2,sorted3,sorted4,sorted5;	
wire signed[3:0]n0,n1,n2,n3,n4,n5;	

wire signed[4:0] k0;
wire signed[4:0] k1;
wire signed[4:0] k2;
wire signed[4:0] k3;
wire signed[4:0] k4;	 
wire signed[4:0] k5;

//==================================================================
// sorting in increasing order sorted0~sorted5
//==================================================================
cmp cmp0 (.A(in_n0 ),.B(in_n1 ),.s(opt[0]),.node0(node00 ),.node1(node01) ); //sort n0,n1
cmp cmp1 (.A(in_n2 ),.B(in_n3 ),.s(opt[0]),.node0(node02 ),.node1(node03) ); //sort n2,n3
cmp cmp2 (.A(in_n4 ),.B(in_n5 ),.s(opt[0]),.node0(node04 ),.node1(node05) ); //sort n4,n5
cmp cmp3 (.A(node00),.B(node02),.s(opt[0]),.node0(node10 ),.node1(node12) ); //sort n0,n2
cmp cmp4 (.A(node10),.B(node04),.s(opt[0]),.node0(sorted0),.node1(node14) ); //sort n0,n4
cmp cmp5 (.A(node01),.B(node05),.s(opt[0]),.node0(node11 ),.node1(node15) ); //sort n1,n5
cmp cmp6 (.A(node03),.B(node15),.s(opt[0]),.node0(node13 ),.node1(sorted5)); //sort n3,n5
cmp cmp7 (.A(node11),.B(node12),.s(opt[0]),.node0(node21 ),.node1(node22) ); //sort n1,n2
cmp cmp8 (.A(node13),.B(node14),.s(opt[0]),.node0(node23 ),.node1(node24) ); //sort n3,n4
cmp cmp9 (.A(node21),.B(node23),.s(opt[0]),.node0(sorted1),.node1(node33) ); //sort n1,n3
cmp cmp10(.A(node22),.B(node24),.s(opt[0]),.node0(node32 ),.node1(sorted4)); //sort n2,n4
cmp cmp11(.A(node32),.B(node33),.s(opt[0]),.node0(sorted2),.node1(sorted3)); //sort n2,n3

//output sort0~sort5

//==================================================================
//cal n0~n5 with opt[1]
//==================================================================
assign n0 = opt[1] ? sorted5 : sorted0; 
assign n1 = opt[1] ? sorted4 : sorted1; 
assign n2 = opt[1] ? sorted3 : sorted2; 
assign n3 = opt[1] ? sorted2 : sorted3; 
assign n4 = opt[1] ? sorted1 : sorted4; 
assign n5 = opt[1] ? sorted0 : sorted5; 

//output n0~n5
//==================================================================
// shifting and moving avg
//==================================================================

assign k0 = {(opt[0]&n0[3]),n0};
assign k1 = {(opt[0]&n1[3]),n1};
assign k2 = {(opt[0]&n2[3]),n2};
assign k3 = {(opt[0]&n3[3]),n3};
assign k4 = {(opt[0]&n4[3]),n4};
assign k5 = {(opt[0]&n5[3]),n5};

wire signed[4:0]div_3_1_result;
wire signed[4:0]div_3_2_result;
wire signed[4:0]div_3_3_result;
wire signed[4:0]div_3_4_result;
wire signed[4:0]div_3_5_result;



wire signed[4:0] neg_k0 = -k0;
	
wire signed[4:0] m0 = opt[2] ?             k0 : 5'b0;

wire signed[6:0]tmp_1 = k1 + k0 * 2;
div_3 div_3_1(.in(tmp_1),.out(div_3_1_result));
wire signed[4:0] m1 = opt[2] ? div_3_1_result : k1 + neg_k0;

wire signed[6:0]tmp_2 = k2 + m1 * 2;
div_3 div_3_2(.in(tmp_2),.out(div_3_2_result));
wire signed[4:0] m2 = opt[2] ? div_3_2_result : k2 + neg_k0;

wire signed[6:0]tmp_3 = k3 + m2 * 2;
div_3 div_3_3(.in(tmp_3),.out(div_3_3_result));
wire signed[4:0] m3 = opt[2] ? div_3_3_result : k3 + neg_k0;

wire signed[6:0]tmp_4 = k4 + m3 * 2;
div_3 div_3_4(.in(tmp_4),.out(div_3_4_result));
wire signed[4:0] m4 = opt[2] ? div_3_4_result : k4 + neg_k0;

wire signed[6:0]tmp_5 = k5 + m4 * 2;
div_3 div_3_5(.in(tmp_5),.out(div_3_5_result));
wire signed[4:0] m5 = opt[2] ? div_3_5_result : k5 + neg_k0;






//result is m0~m5

//==================================================================
// calculate out_n with equ
//==================================================================
wire signed [6:0]add_in1,add_in2;
wire signed [7:0]add_out;


assign add_in1 = equ ? m0 : m3;
assign add_in2 = equ ? -m1 : m4*4;


assign add_out = add_in1 + add_in2;

wire signed[11:0] tmp = m5 * add_out;
wire signed	[10:0]div_result;
div_3_12b div_3_12b_1(tmp,div_result);
assign out_n = (equ&&tmp[11]) ? (-tmp) : (equ ? tmp : div_result);

 



endmodule



module cmp(
	A,
	B,
	s,
	node0,
	node1
);
	input [3:0]A;
	input [3:0]B;
	input s;
	output wire [3:0] node0;
	output wire [3:0] node1;

	wire signed[4:0]e_A = {s&A[3],A};
	wire signed[4:0]e_B = {s&B[3],B};
	
	assign node0 = (e_A<e_B ? A : B);
	assign node1 = (e_A<e_B ? B : A);
	

endmodule