/home/RAID2/COURSE/iclab/iclabta01/umc018/Lef/umc18_6lm.lef